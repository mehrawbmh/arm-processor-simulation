module instruction_Memory(input[31:0] addr, output [31:0] memOut);
    reg [31:0] mem [0:31] ;

    initial begin
        mem[0]=32'b1110_00_1_1101_0_0000_0000_000000010100;
        mem[1]=32'b1110_00_1_1101_0_0000_0001_101000000001;
        mem[2]=32'b1110_00_1_1101_0_0000_0010_000100000011;
        mem[3]=32'b1110_00_0_0100_1_0010_0011_000000000010;
        mem[4]=32'b1110_00_0_0101_0_0000_0100_000000000000;
        mem[5]=32'b1110_00_0_0010_0_0100_0101_000100000100;
        mem[6]=32'b1110_00_0_0110_0_0000_0110_000010100000;
        mem[7]=32'b1110_00_0_1100_0_0101_0111_000101000010;
        mem[8]=32'b1110_00_0_0000_0_0111_1000_000000000011;
        mem[9]=32'b1110_00_0_1111_0_0000_1001_000000000110;
        mem[10]=32'b1110_00_0_0001_0_0100_1010_000000000101;
        mem[11]=32'b1110_00_0_1010_1_1000_0000_000000000110;
        mem[12]=32'b0001_00_0_0100_0_0001_0001_000000000001;
        mem[13]=32'b1110_00_0_1000_1_1001_0000_000000001000;
        mem[14]=32'b0000_00_0_0100_0_0010_0010_000000000010;
        mem[15]=32'b1110_00_1_1101_0_0000_0000_101100000001;
    end

    assign memOut = mem[addr[31:2]];


endmodule