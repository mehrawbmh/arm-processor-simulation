module instruction_Memory(input[31:0] addr, output [31:0] memOut);
    reg [31:0] mem [0:63] ;

    initial begin
        mem[0] = 32'b1110_00_1_1101_0_0000_0000_000000010100;
        mem[1] = 32'b1110_00_1_1101_0_0000_0001_101000000001;
        mem[2] = 32'b1110_00_1_1101_0_0000_0010_000100000011;
        mem[3] = 32'b1110_00_0_0100_1_0010_0011_000000000010;
        mem[4] = 32'b1110_00_0_0101_0_0000_0100_000000000000;
        mem[5] = 32'b1110_00_0_0010_0_0100_0101_000100000100;
        mem[6] = 32'b1110_00_0_0110_0_0000_0110_000010100000;
        mem[7] = 32'b1110_00_0_1100_0_0101_0111_000101000010;
        mem[8] = 32'b1110_00_0_0000_0_0111_1000_000000000011;
        mem[9] = 32'b1110_00_0_1111_0_0000_1001_000000000110;
        mem[10] = 32'b1110_00_0_0001_0_0100_1010_000000000101;
        mem[11] = 32'b1110_00_0_1010_1_1000_0000_000000000110;
        mem[12] = 32'b0001_00_0_0100_0_0001_0001_000000000001;
        mem[13] = 32'b1110_00_0_1000_1_1001_0000_000000001000;
        mem[14] = 32'b0000_00_0_0100_0_0010_0010_000000000010;
        mem[15] = 32'b1110_00_1_1101_0_0000_0000_101100000001;
		mem[16] = 32'b1110_01_0_0100_0_0000_0001_000000000000; //STR		R1 ,[R0],#0	//MEM[1024] = 8192
		mem[17] = 32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR		R11,[R0],#0	//R11 = 8192
		mem[18] = 32'b1110_01_0_0100_0_0000_0010_000000000100; //STR		R2 ,[R0],#4	//MEM[1028] = -1073741824
		mem[19] = 32'b1110_01_0_0100_0_0000_0011_000000001000; //STR		R3 ,[R0],#8	//MEM[1032] = -2147483648
		mem[20] = 32'b1110_01_0_0100_0_0000_0100_000000001101; //STR		R4 ,[R0],#13	//MEM[1036] = 41
		mem[21] = 32'b1110_01_0_0100_0_0000_0101_000000010000; //STR		R5 ,[R0],#16	//MEM[1040] = -123
		mem[22] = 32'b1110_01_0_0100_0_0000_0110_000000010100; //STR		R6 ,[R0],#20	//MEM[1044] = 10
		mem[23] = 32'b1110_01_0_0100_1_0000_1010_000000000100; //LDR		R10,[R0],#4	//R10 = -1073741824
		mem[24] = 32'b1110_01_0_0100_0_0000_0111_000000011000; //STR		R7 ,[R0],#24	//MEM[1048] = -123
		mem[25] = 32'b1110_00_1_1101_0_0000_0001_000000000100; //MOV		R1 ,#4		//R1 = 4
		mem[26] = 32'b1110_00_1_1101_0_0000_0010_000000000000; //MOV		R2 ,#0		//R2 = 0
		mem[27] = 32'b1110_00_1_1101_0_0000_0011_000000000000; //MOV		R3 ,#0		//R3 = 0
		mem[28] = 32'b1110_00_0_0100_0_0000_0100_000100000011; //ADD		R4 ,R0,R3,LSL #2	
		mem[29] = 32'b1110_01_0_0100_1_0100_0101_000000000000; //LDR		R5 ,[R4],#0
		mem[30] = 32'b1110_01_0_0100_1_0100_0110_000000000100; //LDR		R6 ,[R4],#4
		mem[31] = 32'b1110_00_0_1010_1_0101_0000_000000000110; //CMP		R5 ,R6
		mem[32] = 32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGT		R6 ,[R4],#0
		mem[33] = 32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGT		R5 ,[R4],#4
		mem[34] = 32'b1110_00_1_0100_0_0011_0011_000000000001; //ADD		R3 ,R3,#1
		mem[35] = 32'b1110_00_1_1010_1_0011_0000_000000000011; //CMP		R3 ,#3
		mem[36] = 32'b1011_10_1_0_111111111111111111110111      ; //BLT		#-9
		mem[37] = 32'b1110_00_1_0100_0_0010_0010_000000000001; //ADD		R2 ,R2,#1
		mem[38] = 32'b1110_00_0_1010_1_0010_0000_000000000001; //CMP		R2 ,R1
		mem[39] = 32'b1011_10_1_0_111111111111111111110011      ; //BLT		#-13
		mem[40] = 32'b1110_01_0_0100_1_0000_0001_000000000000; //LDR		R1 ,[R0],#0	//R1 = -2147483648
		mem[41] = 32'b1110_01_0_0100_1_0000_0010_000000000100; //LDR		R2 ,[R0],#4	//R2 = -1073741824
		mem[42] = 32'b1110_01_0_0100_1_0000_0011_000000001000; //LDR		R3 ,[R0],#8	//R3 = 41
		mem[43] = 32'b1110_01_0_0100_1_0000_0100_000000001100; //LDR		R4 ,[R0],#12	//R4 = 8192
		mem[44] = 32'b1110_01_0_0100_1_0000_0101_000000010000; //LDR		R5 ,[R0],#16	//R5 = -123
		mem[45] = 32'b1110_01_0_0100_1_0000_0110_000000010100; //LDR		R6 ,[R0],#20	//R6= 10
		mem[46] = 32'b1110_10_1_0_111111111111111111111111      ; //B		#-1
    end

    assign memOut = mem[addr[31:2]];


endmodule